package environment_pkg;

	import uvm_pkg::*;
	
	`include "uvm_macros.svh"

	`include "helpers.svh"

	`include "uart_sequence_item.svh"
	`include "transmitter_sequence_item.svh"
	`include "transmitter_baud_sequence.svh"
	`include "transmitter_reset_sequence.svh"
	`include "transmitter_threshold_sequence.svh"
	`include "transmitter_driver.svh"
	`include "transmitter_input_monitor.svh"
	`include "transmitter_output_monitor.svh"
	`include "transmitter_input_coverage.svh"
	`include "transmitter_output_coverage.svh"
	`include "transmitter_sequencer.svh"
	`include "transmitter_input_agent.svh"
	`include "transmitter_output_agent.svh"
	`include "transmitter_scoreboard.svh"
	`include "transmitter_environment.svh"
   
	
endpackage : environment_pkg
