package test_pkg;

	import uvm_pkg::*;

	`include "uvm_macros.svh"

	import env_pkg::*;

	// Tests
	`include "transmitter_test_base.svh"
	`include "transmitter_basic_test.svh"


endpackage : test_pkg