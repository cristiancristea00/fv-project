class transmitter_sequence_item extends uvm_sequence_item;

    `uvm_object_utils(transmitter_sequence_item)

    function new(string name = "transmitter_sequence_item");
        super.new(name);
    endfunction


    rand  bit               write_enable;
    randc bit [7:0]         data;
    rand  bit [5:0]         buffer_full_threshold;
    rand  baudrate_select_t baudrate_select;


    constraint buffer_full_threshold_constraint {
        buffer_full_threshold == 32;
    }

    constraint baudrate_select_constraint {
        baudrate_select == BAUD_CLK16;
    }

    constraint write_enable_constraint {
        write_enable == 1;
    }


    function void kill();
        write_enable          = 0;
        data                  = 0;
        buffer_full_threshold = 32;
        baudrate_select       = BAUD_CLK16;
    endfunction: kill


    virtual function void do_print(uvm_printer printer);
        printer.print_int("baudrate_select", baudrate_select, $bits(baudrate_select), UVM_DEC, ".", "dec");
        printer.print_int("buffer_full_threshold", buffer_full_threshold, $bits(buffer_full_threshold), UVM_DEC, ".", "dec");
        printer.print_string("data", get_data_str());
        printer.print_string("uart_data", get_uart_data_str());
        printer.print_string("write_enable", write_enable ? "True" : "False");
    endfunction: do_print


    function string get_data_str();
        string data_str = $sformatf("%h", data);

        return $sformatf("0x%s", data_str.toupper());
    endfunction: get_data_str


    function string get_uart_data_str();
        return $sformatf("%b", get_uart_data());
    endfunction: get_uart_data_str


    function bit[8:0] get_uart_data();
        return {data[0], data[1], data[2], data[3], data[4], data[5], data[6], data[7], ^data};
    endfunction: get_uart_data


endclass: transmitter_sequence_item
