

class uart_seq_item extends uvm_sequence_item;
   `uvm_object_utils(uart_seq_item)
   
   
   function new(string name= "uart_seq_item");
      super.new(name);
   endfunction



endclass: uart_sequence_item
