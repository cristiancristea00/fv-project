
interface sys_itf();


 
// Write initial reset here 
    initial begin

    end

//Initialise required signals with 0 here
    initial begin
    
    end
 
// Complete this task in order to implement the reset task 
    task drive_reset(int len);

    endtask: drive_reset
   
endinterface
