package tests_pkg;

	import uvm_pkg::*;

	`include "uvm_macros.svh"

	import environment_pkg::*;

	// Tests
	`include "transmitter_test_base.svh"
	`include "transmitter_basic_test.svh"


endpackage : tests_pkg