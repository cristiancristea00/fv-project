package tests_pkg;

	import uvm_pkg::*;

	`include "uvm_macros.svh"

	import environment_pkg::*;

	`include "transmitter_base_test.svh"
	`include "transmitter_basic_test.svh"


endpackage : tests_pkg