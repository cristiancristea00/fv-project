package env_pkg;

	import uvm_pkg::*;
	
	`include "uvm_macros.svh"
   
endpackage : env_pkg
