
`include "uvm_macros.svh"


 import  uvm_pkg::*; 

  
module uart_transmitter_tb();


logic rst_n_s;


// Generate clock signal here or as a separate module
initial begin

end


 
// Connect all the required signals below


// Upload the interface to the UVM_CONFIG_DB here
initial begin
	
	run_test("");
end

endmodule
